module hello_world;
initial
begin
	$display("hello_world");
	#10 $finish;
end

endmodule